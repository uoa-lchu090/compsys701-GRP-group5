package ram_constants is
	
	constant ram_addr_width: integer := 10;
	constant ram_data_width: integer := 16;
	
	constant rom_addr_width: integer := 10;
	constant rom_data_width: integer := 32;

end ram_constants;